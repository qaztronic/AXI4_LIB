// --------------------------------------------------------------------
// Copyright 2024 qaztronic
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
// Licensed under the Solderpad Hardware License v 2.1 (the “License”);
// you may not use this file except in compliance with the License, or,
// at your option, the Apache License version 2.0. You may obtain a copy
// of the License at
//
// https://solderpad.org/licenses/SHL-2.1/
//
// Unless required by applicable law or agreed to in writing, any work
// distributed under the License is distributed on an “AS IS” BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or
// implied. See the License for the specific language governing
// permissions and limitations under the License.
// --------------------------------------------------------------------

module clocks_ratio #(N=2, W=16)
( input              clk
, input              reset
, input              trigger
, input              clk_in[N]
, output reg [W-1:0] count [N]
);
  // --------------------------------------------------------------------
  wire trigger_z[N];
  wire rise_edge[N];
  wire fall_edge[N];

  generate
    for(genvar j = 0; j < N; j = j + 1)
    begin: sync
      half_synchronizer
        half_synchronizer_i
        ( .in       (trigger     )
        , .out_clk  (clk_in [j]  )
        , .out      (trigger_z[j])
        , .rise_edge(rise_edge[j])
        , .fall_edge(fall_edge[j])
        );
    end
  endgenerate

  // --------------------------------------------------------------------
  wire [N-1:0] overflow;
  wire any_overflow = |overflow;

  generate
    for(genvar j = 0; j < N; j = j + 1)
    begin: counter
      assign overflow[j] = &count[j];

      always_ff @(posedge clk_in[j])
        if(reset | rise_edge[j])
          count[j] = 0;
        else if(~overflow[j] & ~any_overflow)
          count[j] = count[j] + 1;
    end
  endgenerate

// --------------------------------------------------------------------
endmodule
