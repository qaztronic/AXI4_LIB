// -----------------------------------------------------------------------------
// Copyright qaztronic    |    SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
// Licensed under the Solderpad Hardware License v 2.1 (the "License"); you may
// not use this file except in compliance with the License, or, at your option,
// the Apache License version 2.0. You may obtain a copy of the License at
// https://solderpad.org/licenses/SHL-2.1/
//
// Unless required by applicable law, any work distributed under the License is
// distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY
// KIND, either express or implied. See the License for the specific language
// governing permissions and limitations under the License.
// -----------------------------------------------------------------------------

// --------------------------------------------------------------------
package axi4_lite_pkg;
  // --------------------------------------------------------------------
  typedef struct packed {
    int A;
    int N;
    int I;
    int USE_STRB;
    int USE_PROT;
    int USE_MOD_PORT;
  } axi4_lite_cfg_t;

// --------------------------------------------------------------------
endpackage
