// --------------------------------------------------------------------
// Copyright 2024 qaztronic
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
// Licensed under the Solderpad Hardware License v 2.1 (the “License”);
// you may not use this file except in compliance with the License, or,
// at your option, the Apache License version 2.0. You may obtain a copy
// of the License at
//
// https://solderpad.org/licenses/SHL-2.1/
//
// Unless required by applicable law or agreed to in writing, any work
// distributed under the License is distributed on an “AS IS” BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or
// implied. See the License for the specific language governing
// permissions and limitations under the License.
// --------------------------------------------------------------------

module half_synchronizer #(W=3)
( input  in
, input  out_clk
, output out
, output rise_edge
, output fall_edge
);
  // --------------------------------------------------------------------
  reg [W:0] out_r;
  assign out = out_r[1];
  assign rise_edge = ~out_r[0] &  out_r[1];
  assign fall_edge =  out_r[0] & ~out_r[1];

  always_ff @(posedge out_clk)
    out_r <= {in, out_r[W:1]};

// --------------------------------------------------------------------
endmodule
